*Simulation of CMOS inverter
M1 2 1 0 0 MOSN W=5U L=1.0U
M2 2 1 3 3 MOSP W=5U L=1.0U
VIN 1 0 DC 5V PULSE (0 5V 0 1NS 1NS 20US 40US)
VDD 3 0 DC 5.0
.MODEL MOSN NMOS VTO=0.7 KP=110U GAMMA=0.4 LAMBDA=0.04 PHI=0.7
.MODEL MOSP PMOS VTO=-0.7 KP=50U GAMMA=0.57 LAMBDA=0.05 PHI=0.8
.TRAN 1US 100US
.OP
.PRINT TRAN V(2) V(1)
.PROBE
.END
