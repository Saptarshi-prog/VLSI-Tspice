*CMOS inverter with a load capacitance of 50fF
M1 2 1 0 0 MOSN W=5U L=1.0U
M2 2 1 3 3 MOSP W=12.5U L=1.0U
VIN 1 0 DC 5V PULSE(0 5V 0 0.1PS 0.1PS 200PS 400PS)
VDD 3 0 DC 5.0
C 2 0 50fF
.MODEL MOSN NMOS VTO=0.7 KP=110U GAMMA=0.4 LAMBDA=0.04 PHI=0.7
.MODEL MOSP PMOS VTO=-0.7 KP=44U GAMMA=0.57 LAMBDA=0.05 PHI=0.8
.TRAN 1PS 800PS
.OP
.PRINT TRAN V(2) V(1)
.PROBE
.END