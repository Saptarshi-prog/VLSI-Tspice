M1 1 3 4 0 MOSN W=0.8U L=0.2U
M2 4 2 1 5 MOSP W=0.4U L=0.2U
M3 4 2 10 0 MOSN W=0.8U L=0.2U
M4 10 3 4 5 MOSP W=0.4U L=0.2U

M5 9 4 0 0 MOSN W=0.8U L=0.2U
M6 9 4 5 5 MOSP W=0.4U L=0.2U
M7 10 9 0 0 MOSN W=0.8U L=0.2U
M8 10 9 5 5 MOSP W=0.4U L=0.2U

C 10 0 10fF

*Control SigNl
VC1 3 0 DC 5V PULSE(0 5V 0 0 0 100PS 200PS)
VC2 2 0 DC 5V PULSE(5V 0 0 0 0 100PS 200PS)

*Input Signal
VIN 1 0 DC 5V PULSE(0 5V 0 0 0 175PS 400PS)

VDD 5 0 DC 5.0
.MODEL MOSN NMOS VTO=0.5 KP=270U GAMMA=0.3 LAMBDA=0.04 PHI=0.84
.MODEL MOSP PMOS VTO=-0.5 KP=70U GAMMA=0.3 LAMBDA=0.05 PHI=0.84
.TRAN 0.5PS 1200PS
.OP
.PRINT TRAN v(10) 
.PROBE
.END
