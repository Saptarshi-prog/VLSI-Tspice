*Simulation of CMOS NAND Gate
M1 5 1 0 0 MOSN W=5U L=1.0U
M2 3 2 5 5 MOSN W=5U L=1.0U
M3 3 2 4 4 MOSP W=5U L=1.0U
M4 3 1 4 4 MOSP W=5U L=1.0U
VA 2 0 DC 5V PULSE(0 5V 0 1NS 1NS 20US 40US)
VB 1 0 DC 5V PULSE(0 5V 0 1NS 1NS 30US 40US)
VDD 4 0 DC 5.0
.MODEL MOSN NMOS VTO=0.7 KP=110U GAMMA=0.4 LAMBDA=0.04 PHI=0.7
.MODEL MOSP PMOS VTO=-0.7 KP=50U GAMMA=0.57 LAMBDA=0.05 PHI=0.8
.TRAN 1US 150US
.OP
.PRINT TRAN V(3) V(2) V(1)
.PROBE
.END
